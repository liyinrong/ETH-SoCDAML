`include "tmicro-classes.sv"
`define NUM_INSTRUCTIONS 80

class nml_program;
    rand tmicro$tmicro moves[20];
    rand tmicro$tmicro ariths[`NUM_INSTRUCTIONS];
    rand tmicro$tmicro halt;
    function new();
        foreach (moves[i]) moves[i] = new();
        foreach (ariths[i]) ariths[i] = new();
        halt = new();
    endfunction
    function print(int out_file);
        foreach (moves[i])
          $fdisplay(out_file, moves[i].get_bits_and_syntax());
        foreach (ariths[i])
          $fdisplay(out_file, ariths[i].get_bits_and_syntax());
        $fdisplay(out_file, halt.get_bits_and_syntax());
    endfunction
    constraint c {
        // First move some random values into registers
        foreach (moves[i])
            (moves[i].sub == tmicro$tmicro::S$move_instr &&
             moves[i].R$move_instr.sub == tmicro$move_instr::S$mvi_wreg_word &&
             moves[i].R$move_instr.R$mvi_wreg_word.P$rr.sub == tmicro$wreg::S$r_reg);
        // Now perform some random additions
        foreach (ariths[i])
            (ariths[i].sub == tmicro$tmicro::S$alu_instr &&
             ariths[i].R$alu_instr.sub == tmicro$alu_instr::S$alu_rrr &&
             ariths[i].R$alu_instr.R$alu_rrr.P$op.val == tmicro$alu_op$0::E$add &&
             ariths[i].R$alu_instr.R$alu_rrr.P$t.P$r.val inside {[0:3]});
        // Finally, a halt instruction
        (halt.sub == tmicro$tmicro::S$control_instr &&
         halt.R$control_instr.sub == tmicro$control_instr::S$halt);
    }
endclass;


program main;
   initial begin
       nml_program prog;
       string filename = "risk_tmicro_sv.ras";
       int out_file = $fopen(filename);
       $display("Generating instructions in \"%s\"", filename);
       $fdisplay (out_file, "// Generated by SystemVerilog by Risk");
       $fdisplay (out_file, "");
       $fdisplay (out_file, ".text_segment PM 0");
       prog = new();
       prog.randomize();
       prog.print(out_file);
       $fclose(out_file);
   end
endprogram
